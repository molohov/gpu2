module gpu (
    input polygon,
    output framebuffer
);

// insert gpu code here
assign framebuffer = polygon;

endmodule
